
library ieee;
use ieee.std_logic_1164.all;

entity CPU is
end entity CPU;
